`ifndef ENUMS

//ALU Enums
parameter e_ALU_noop = 0;
parameter e_ALU_add = 1;
parameter ALU_OP_W = 1;

`define ENUMS
`endif

// This file is dynamically generated to just point to the file where our binary is stored
// the include path should be relative to the location of this file
`include "../output/binary.vh"